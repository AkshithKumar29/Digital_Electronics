`timescale 1ns/1ps
module tb_full_subtractor_using_half_subtractor;
    reg A, B, Bin;
    wire D, Bout; 
    full_subtractor_using_half_subtractor uut(.A(A), .B(B), .Bin(Bin), .D(D), .Bout(Bout));
    initial begin
        $dumpfile("full_subtractor_using_half_subtractor.vcd");
        $dumpvars(0, tb_full_subtractor_using_half_subtractor);
        $monitor("Time = %0t, A = %b, B = %b, Bin = %b -> D = %b, Bout = %b", $time,A,B,Bin,D,Bout);
        A = 0; B = 0; Bin = 0; #10;
        A = 0; B = 0; Bin = 1; #10;
        A = 0; B = 1; Bin = 0; #10;
        A = 0; B = 1; Bin = 1; #10;
        A = 1; B = 0; Bin = 0; #10;
        A = 1; B = 0; Bin = 1; #10;
        A = 1; B = 1; Bin = 0; #10;
        A = 1; B = 1; Bin = 1; #10;
    end
endmodule