module full_adder(

);
endmodule